// Bit and register definitions for test_control module
//
// 13-Feb-2019 DFN Initial version to improve documentation

`define USE_FAKE_ADDR 0
 `define USE_FAKE_PPS_BIT 0
 `define USE_FAKE_SHWR_BIT 1
 `define USE_FAKE_MUON_BIT 2
 `define USE_FAKE_RD_BIT 3
 `define USE_FAKE_RDCLK_BIT 4
 `define DISABLE_TRIG_OUT_BIT 5

 `define FAKE_MODE_ADDR 1
