`ifndef _TRIGGER_OPTIONS
  `define _TRIGGER_OPTIONS
  `define COMPILE_DATE 'h10050319
`endif
