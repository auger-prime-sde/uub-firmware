`ifndef _RD_IFC_OPTIONS
  `define _RD_IFC_OPTIONS
  `define RD_IFC_COMPILE_DATE 'h19151120
`endif
