`ifndef _TRIGGER_OPTIONS
  `define _TRIGGER_OPTIONS
  `define COMPILE_DATE 'h18081119
`endif
