// Header file for module to configure the digital interfaces
//
// 24-Mar-2019 DFN Initial version

// Digital Interface register assignments
`define DIG_IFC_CONTROL_ADDR 0
`define DIG_IFC_INPUT_ADDR 1
`define DIG_IFC_OUTPUT_ADDR 2
`define DIG_IFC_ID_ADDR 3
