`ifndef _TRIGGER_OPTIONS
  `define _TRIGGER_OPTIONS
  `define COMPILE_DATE 'h20090719
`endif
